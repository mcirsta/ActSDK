cdl_package CYGPKG_NORMAL_CONFIG {
	display			"������Ϣ����"
	define_header 	tools.gn
	description		"configuration item for fw tools"
	
	define_proc {
		puts $::cdl_header "#include \"tools_inner.h\""
		puts $::cdl_header ""
	}

	cdl_component USB_CFG {
		display "USB �������"
		flavor none
		no_define
		description "����USB��ص�����"
		
		define_proc {
			puts $::cdl_header ""
			puts $::cdl_header "/*USB�������*/"
		}
		
		cdl_option PID {
			display "PID"
			flavor data
			no_define
			default_value {"PID=0x1101"}
			define ADDCONFIG
			
			define_proc {
				puts $::cdl_header "/*end of PID*/"
				puts $::cdl_header ""
			}
		}
		
		
		cdl_option VID {
			display "VID"
			flavor data
			no_define
			default_value {"VID=0x10D6"}
			define ADDCONFIG
			
			define_proc {
				puts $::cdl_header "/*end of VID*/"
				puts $::cdl_header ""
			}
		}
		
		cdl_option USBATTRI {
			display "USB ����"
			flavor data
			default_value {"USBATTRI_8=\"GENERIC\""}
			no_define
			define 	ADDCONFIG
			description "
				����USB���ԣ�ע�⣺valueֵ���ַ���󳤶�Ϊ8.
				"
			define_proc {
				puts $::cdl_header ""
			}
		}
		
		cdl_option USBIDENTIFICATION {
			display "USB ID"
			flavor data
			default_value {"USBIDENTIFICATION_16=\"USB DISK DEVICE\""}
			no_define
			define ADDCONFIG
			description "����USB ID��ע�⣺VALUEֵ���ַ���󳤶�Ϊ16"
			define_proc {
				puts $::cdl_header ""
			}
		}
		
		cdl_option USBPRODUCTVER {
			display "USB��Ʒ�汾"
			flavor data
			default_value {"USBPRODUCTVER_4=\"1.00\""}
			no_define
			define ADDCONFIG
			description "����USB��Ʒ�汾�ţ�ע�⣺VALUEֵ���ַ���󳤶�Ϊ4"
			define_proc {
				puts $::cdl_header ""
			}
		}
		
		cdl_option USBDESCRIPSTR {
			display "USB������Ϣ"
			flavor data
			default_value {"USBDESCRIPSTR_23=\"USB MASS STORAGE CLASS\""}
			no_define
			define ADDCONFIG
			description "USB������Ϣ��ע�⣺VALUEֵ���ַ���󳤶�Ϊ23"
			define_proc {
				puts $::cdl_header ""
			}
		}
		
		cdl_option USBSERIAL {
			display "U���Ƿ��ϱ���Ʒ���к�"
			flavor data
			default_value {"UdiskSerialNumFlag=1"}
			no_define
			define ADDCONFIG
			description "U�����Ƿ��ϱ���Ʒ���кţ�0-no��1-yes��"
			define_proc {
				puts $::cdl_header ""
			}
		}
	}
	
	cdl_component MTP_CFG {
		display "MTP �������"
		flavor none
		no_define
		description "MTP�������"
	
		cdl_option MTPPID {
			display "MTPPID"
			flavor data
			no_define
			default_value {"MTPPID=0x2300"}
			define ADDCONFIG
			
			define_proc {
				puts $::cdl_header "/*end of MTPPID*/"
				puts $::cdl_header ""
			}
		}
		
		
		cdl_option MTPVID {
			display "MTPVID"
			flavor data
			no_define
			default_value {"MTPVID=0x10D6"}
			define ADDCONFIG
			
			define_proc {
				puts $::cdl_header "/*end of MTPVID*/"
				puts $::cdl_header ""
			
			}
		}
		
		cdl_option MTPMFTINFO {
			display "MTPMFTINFO����"
			flavor data
			default_value {"MTPMFTINFO=\"Actions Semiconductor Co., Ltd.\""}
			no_define
			define ADDCONFIG
			description "MTPMFTINFO����,ע�⣺VALUEֵ���ַ���󳤶�Ϊ32"
			
			define_proc {
				puts $::cdl_header ""
			}
		}
		
		cdl_option MTPPRODUCTINFO {
			display "MTPPRODUCTINFO����"
			flavor data
			default_value {"MTPPRODUCTINFO=\"Actions Mtp Device 000001\""}
			no_define
			define ADDCONFIG
			description "MTPPRODUCTINFO����,ע�⣺VALUEֵ���ַ���󳤶�Ϊ32"
			
			define_proc {
				puts $::cdl_header ""
			}
		}
		
		cdl_option MTPPRODUCTVER {
			display "MTPPRODUCTVER����"
			flavor data
			default_value {"MTPPRODUCTVER=\"V1.00.3333\""}
			no_define
			define ADDCONFIG
			description "MTPPRODUCTVER����,ע�⣺VALUEֵ���ַ���󳤶�Ϊ16"
			
			define_proc {
				puts $::cdl_header ""
			}
		}
	}

	cdl_component NandFlashCE_CFG {
		display "NandFlashCE ����"
		no_define
		description "����4CE�������Ƭѡ��Ϣ"
		
		cdl_option NandflashCE_TYPE {
			display "NandFlash CE��������"
			flavor data
			default_value 1
			legal_values {1 2}
			no_define
			description "1��gpio��ʽ��2��MUX��ʽ"
		}
		
		cdl_option NandflashCE_RESERVE {
			display "NandFlash CE��������"
			flavor data
			default_value 0
			no_define
			description "��ʱ��������"
		}
		
		cdl_option NandflashCE_CE3 {
			display "Nandflash CE3ʵ�ַ�ʽ"
			flavor data
			no_define
			description "0��31ΪgpioA��id��32��63ΪgpioB�Ķ�Ӧid"
		}
		
		cdl_option NandflashCE_CE4 {
			display "Nandflash CE4ʵ�ַ�ʽ"
			flavor data
			no_define
			description "0��31ΪgpioA��id��32��63ΪgpioB�Ķ�Ӧid"
		}
		
		
		cdl_option NandflashCE_CFG {
			display "NandFlash ����"
			flavor data
			calculated { (NandflashCE_TYPE<<24) + (NandflashCE_RESERVE<<16)+ (NandflashCE_CE3<<8) + NandflashCE_CE4 }
			no_define
			define ADDAFINFO_VALUE
			description "dNandflashCE ����"
			
			define_proc {
				puts $::cdl_header "#define ADDAFINFO_OFFSET 0x180"
				puts $::cdl_header "#define ADDAFINFO_LEN 0x4"
				puts $::cdl_header "/*end of NandflashCE_CFG*/"
				puts $::cdl_header ""
			}
		}
	}
	
	cdl_option RTC_SOURCE {
		display 	"RTC ʱ��Դ����"
		flavor data
		default_value 0
		legal_values {0 1}
		description "RTC ʱ��Դ���ã� \n
			0�� �ⲿʱ��Դ	\n
			1�� �ڲ�ʱ��Դ	\n"
		no_define
		define ADDFMINFO_VALUE
		
		define_proc {
			puts $::cdl_header "#define ADDFMINFO_OFFSET 0x42"
			puts $::cdl_header "#define ADDFMINFO_LEN 0x4"
			puts $::cdl_header "/*end of RTC_SOURCE*/"
			puts $::cdl_header ""
		}
	}

	
	cdl_option VER {
		display "���̹̼��汾��"
		flavor data
		no_define
		default_value {"VER=\"13.00.10.1017.20080515\""}
		define ADDCONFIG
		
		define_proc {
			puts $::cdl_header "/*end of VER*/"
			puts $::cdl_header ""
		}
	}

	cdl_option SCODE_CAP {
		display "ϵͳ��������С(��λ������)"
		flavor data
		default_value 1
		no_define
		define ADDAFINFO_VALUE
		
		define_proc {
			puts $::cdl_header "#define ADDAFINFO_OFFSET 0x200"
			puts $::cdl_header "#define ADDAFINFO_LEN 0x4"
			puts $::cdl_header "/*end of SCODE_CAP*/"
			puts $::cdl_header ""
		}
	}
	
	
	cdl_option SCODE_CAP_BAK {
		display "ϵͳ���뱸������С(��λ������)"
		flavor data
		default_value 1
		no_define
		define ADDAFINFO_VALUE
		
		define_proc {
			puts $::cdl_header "#define ADDAFINFO_OFFSET 0x204"
			puts $::cdl_header "#define ADDAFINFO_LEN 0x4"
			puts $::cdl_header "/*end of SCODE_CAP_BAK*/"
			puts $::cdl_header ""
		}
	}
	
	
	cdl_option CFG_DEFAULTDATE {
		display "ȱʡ��������"
		flavor data
		default_value {"DATE=\"2000-01-01\""} 
		no_define
		define ADDCONFIG
		define_proc {
			puts $::cdl_header ""
		}
	}
	
	
	cdl_option CFG_DEFAULTTIME {
		display "ȱʡʱ������"
		flavor data
		default_value {"TIME=\"00:00\""} 
		no_define
		define ADDCONFIG
		define_proc {
			puts $::cdl_header ""
		}
	}
	
	
	cdl_option TIME_FORMAT {
		display "ʱ����ʽ����"
		flavor data
		default_value {"TIME_FORMAT=24"} 
		no_define
		define ADDCONFIG
		description "ʱ����ʽ��12/24"
		
		define_proc {
			puts $::cdl_header ""
		}
	}
	
	cdl_option  BACKLIGHT_BRIGHT {
		display "����ѡ��"
		flavor data
		default_value {"BACKLIGHT_BRIGHTNESS=3"} 
		no_define
		define ADDCONFIG
		description "���ȵȼ���1~5"
		
		define_proc {
			puts $::cdl_header ""
		}
	}
	
	
	cdl_option  BACKLIGHT_DURATION {
		display "��������ʱ������"
		flavor data
		default_value {"BACKLIGHT_DURATION=0"} 
		no_define
		define ADDCONFIG
		description "0~60��,����5��"
		
		define_proc {
			puts $::cdl_header ""
		}
	}
		
	cdl_option  IDLE_TIME {
		display "StandBy��ʱ"
		flavor data
		default_value {"IDLE_TIME=0"} 
		no_define
		define ADDCONFIG
		description "0~60��"
		
		define_proc {
			puts $::cdl_header ""
		}
	}
	
	cdl_option  SLEEP_TIME {
		display "˯��ʱ������"
		flavor data
		default_value {"SLEEP_TIME=0"} 
		no_define
		define ADDCONFIG
		description "0~120����"
		
		define_proc {
			puts $::cdl_header ""
		}
	}
	
	cdl_option  LANG_ID {
		display "������������"
		flavor data
		default_value {"LANG_ID=2"} 
		no_define
		define ADDCONFIG
		description "��������, Ӣ��:0, Reserved:1, ����:2 ����:3"
		
		define_proc {
			puts $::cdl_header ""
		}
	}
	
	cdl_option  VOICE_VOLUM {
		display "�����ȼ�����"
		flavor data
		default_value {"VOICE_VOLUM=15"} 
		no_define
		define ADDCONFIG
		description "����, 0~31"
		
		define_proc {
			puts $::cdl_header ""
		}
	}
	
}