cdl_package CYGPKG_APPS_CONFIG {
	display			"Ӧ�ò�������"
	define_header 	tools.gn
	description		"apps configuration item"
	
	cdl_component PHOTO_CFG {
		display "PHOTO �������"
		flavor none
		no_define
		description "PHOTO���ѡ�������"
		
		define_proc {
			puts $::cdl_header ""
			puts $::cdl_header "/*PHOTO�������*/"
		}
		
		cdl_option photo_playmode {
			display "play mode"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1"}
			define -format "photo_playmode=%d" ADDCONFIG
			description "ͼƬ�����ʽ��0-�ֶ������1-�Զ����"
		}
		
		cdl_option photo_browsemode {
			display "browse mode"
			flavor data
			no_define
			default_value {"1"}
			legal_values {"0" "1"}
			define -format "photo_browsemode=%d" ADDCONFIG
			description "�ļ������ʽ��0-�ļ��������1-����ͼ���"
		}
		
		cdl_option photo_slide_effect_mode {
			display "slide effect mode"
			flavor data
			no_define
			default_value {"7"}
			legal_values {"0" "1" "2" "3" "4" "5" "6" "7"}
			define -format "photo_slide_effect_mode=%d" ADDCONFIG
			description "ͼƬ��Ч��ʽ��0-none;1-fade;2-check;3-cut;4-erase;5-louver;6-randomline; 7-random"
		}
		
		cdl_option photo_delaytime {
			display "delay time"
			flavor data
			no_define
			default_value {"2"}
			legal_values {"1" "2" "3" "4" "5" "6" "7" "8" "9" "10"}
			define -format "photo_delaytime=%d" ADDCONFIG
			description "�õ�Ƭ���ż��ʱ�䣺1s~10s"
		}
		
		cdl_option photo_tvout {
			display "photo tvout"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1"}
			define -format "photo_tvout=%d" ADDCONFIG
			description "tvout�����0-off; 1-on"
		}
		
		cdl_option photo_nowplayindex {
			display "nowplay index"
			flavor data
			no_define
			default_value {"0"}
			define -format "photo_nowplayindex=%d" ADDCONFIG
			description "��ǰ����ͼƬ��ƫ��"
		}
		
		cdl_option photo_nowplayname {
			display "nowplay name"
			flavor data
			no_define
			default_value {"a"}
			define -format "photo_nowplayname=\"%s\"" ADDCONFIG
			description "��ǰ����ͼƬ������"
		}
		
		cdl_option photo_nowplaypath {
			display "nowplay path"
			flavor data
			no_define
			default_value {"a"}
			define -format "photo_nowplaypath=\"%s\"" ADDCONFIG
			description "��ǰ����ͼƬ��·��"
		}

	}
		
	cdl_component FM_CFG {
		display "FM �������"
		flavor none
		no_define
		description "FM���ѡ�������"
		
		define_proc {
			puts $::cdl_header ""
			puts $::cdl_header "/*FM�������*/"
		}
		
		cdl_option fm_frequency {
			display "Frequency"
			flavor data
			no_define
			default_value {"87000"}
			define -format "fm_frequency=%d" ADDCONFIG
			description "��ǰ����Ƶ��"
		}
		
		cdl_option fm_band {
			display "Band"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1"}
			define -format "fm_band=%d" ADDCONFIG
			description "�������ã�0- USA Band; 1-JAPAN Band"
		}
		
		cdl_option fm_stereo_mode {
			display "stereo mode"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1"}
			define -format "fm_stereo_mode=%d" ADDCONFIG
			description "������0-mono track;1-stereo track"
		}
		
		cdl_option fm_intensity {
			display "intensity"
			flavor data
			no_define
			default_value {"6"}
			define -format "fm_intensity=%d" ADDCONFIG
			description "������"
		}
		
		cdl_option fm_record_fidelity {
			display "record fidelity"
			flavor data
			no_define
			default_value {"1"}
			legal_values {"0" "1" "2"}
			define -format "fm_record_fidelity=%d" ADDCONFIG
			description "ǿ��:0-low;1-medium;2-hight"
		}
		
		cdl_option fm_record_gain {
			display "record gain"
			flavor data
			no_define
			default_value {"4"}
			legal_values {"1" "2" "3" "4" "5" "6" "7"}
			define -format "fm_record_gain=%d" ADDCONFIG
			description "����:0~7"
		}
			
	}
	
	cdl_component CAMERA_CFG {
		display "CAMERA �������"
		flavor none
		no_define
		description "CAMERA���ѡ�������"
		
		define_proc {
			puts $::cdl_header ""
			puts $::cdl_header "/*CAMERA�������*/"
		}
		
	    cdl_component DC_CFG {
		    display "DC �������"
		    flavor none
		    no_define
		    description "DC���ѡ�������"
		
		    define_proc {
			    puts $::cdl_header ""
			    puts $::cdl_header "/*DC�������*/"
		    }
		
		    cdl_option dc_whitebalance {
			    display "white balance"
			    flavor data
			    no_define
			    default_value {"1"}
			    legal_values {"1" "2" "3" "4" "5"}
			    define -format "dc_whitebalance=%d" ADDCONFIG
			    description "��ƽ��: 1-Auto; 2-Fine; 3-Cloudy; 4-Filament Lamp; 5-Fluorescent Lamp"
		    }
		
		    cdl_option dc_brightness {
			    display "brightness"
			    flavor data
			    no_define
			    default_value {"1"}
			    legal_values {"-3" "-2" "-1" "0" "1" "2" "3" }
			    define -format "dc_brightness=%d" ADDCONFIG
			    description "������: -3~3"
		    }
		
		    cdl_option dc_exposure_mode {
			    display "exposure mode"
			    flavor data
			    no_define
			    default_value {"1"}
			    legal_values {"1" "2" "3"}
			    define -format "dc_exposure_mode=%d" ADDCONFIG
			    description "�ع�ģʽ: 1- Auto; 2-Indoor; 3-Outdoor"
		    }
		
		    cdl_option dc_flashlamp {
			    display "flashlamp"
			    flavor data
			    no_define
			    default_value {"1"}
			    legal_values {"1" "2" "3"}
			    define -format "dc_flashlamp=%d" ADDCONFIG
			    description "�����: 1-Auto; 2-ON; 3-OFF"
		    }
		
		    cdl_option dc_face_identify {
			    display "face identify"
			    flavor data
			    no_define
			    default_value {"1"}
			    legal_values {"1" "2"}
			    define -format "dc_face_identify=%d" ADDCONFIG
			    description "�������: 1-OFF; 2-ON"
		    }
		
		    cdl_option dc_stickerphoto {
		    	display "sticker photo"
		    	flavor data
			    no_define
			    default_value {"1"}
			    legal_values {"1" "2" "3" "4"}
			    define -format "dc_stickerphoto=%d" ADDCONFIG
			    description "��ͷ��: 1-OFF; 2-Photo1; 3-Photo2; 4-Photo3"
		    }
		
		    cdl_option dc_specialeffect {
		    	display "special effect"
		    	flavor data
		    	no_define
		    	default_value {"1"}
		    	legal_values {"1" "2" "3" "4"}
			    define -format "dc_specialeffect=%d" ADDCONFIG
		    	description "��Ч: 1-OFF; 2-Black & White; 3-Sepia; 4-Negative"
		    }
		
		    cdl_option dc_savepath {
		    	display "save path"
		    	flavor data
			    no_define
			    default_value {" "}
			    define -format "dc_savepath=\"%s\"" ADDCONFIG
			    description "����·��"
		    }
		
		    cdl_option dc_resolution {
			    display "resolution"
			    flavor data
			    no_define
			    default_value {"1"}
			    legal_values {"1" "2" "3" "4" "5" "6" "7" "8" "9" "10" "11" "12"}
			    define -format "dc_resolution=%d" ADDCONFIG
			    description "�ֱ���:1.4672x3504; 2.4416x3312; 3.3840x2880; 4.3264x2448; 5.2816x2112; 6.2560x1920; 7.2400x1800; 8.2048x1536; 9.1600x1200; 10.1280x960; 11.1024x768; 12.640x480"
		    }
		
		    cdl_option dc_selftimer {
		    	display "self timer"
		    	flavor data
		    	no_define
		    	default_value {"1"}
		    	legal_values {"1" "2" "3" "4" "5"}
			    define -format "dc_selftimer=%d" ADDCONFIG
		    	description "��ʱ����:1-OFF; 2-5 Sec; 3-10 Sec; 4-15 Sec; 5-20 Sec"
		    }
		
		    cdl_option dc_contshooting {
		    	display "contshooting"
		    	flavor data
		    	no_define
		    	default_value {"1"}
		    	legal_values {"1" "2" "3" "4" "5"}
			    define -format "dc_contshooting=%d" ADDCONFIG
		    	description "��ʱ����:1-OFF; 2-5 Sec; 3-10 Sec; 4-15 Sec; 5-20 Sec"
		    }
		
		    cdl_option dc_shutter_sound {
		    	display "shutter sound"
		    	flavor data
		    	no_define
		    	default_value {"1"}
		    	legal_values {"1" "2" "3" "4"}
			    define -format "dc_shutter_sound=%d" ADDCONFIG
		    	description "��������:1-OFF; 2-Sound1; 3-Sound2; 4-Sound3"
		    }
		
		    cdl_option dc_dater {
		    	display "dater"
		    	flavor data
		    	no_define
		    	default_value {"1"}
		    	legal_values {"1" "2" "3"}
			    define -format "dc_dater=%d" ADDCONFIG
		    	description "���ڱ��:1-OFF; 2-Date; 3-Date & Time"
		    }

	    }
	    cdl_component DV_CFG {
		    display "DV �������"
		    flavor none
		    no_define
		    description "DV���ѡ�������"
		
		    define_proc {
			    puts $::cdl_header ""
			    puts $::cdl_header "/*DV�������*/"
		    }
		    
		    cdl_option dv_whitebalance {
			    display "white balance"
			    flavor data
			    no_define
			    default_value {"1"}
			    legal_values {"1" "2" "3" "4" "5"}
			    define -format "dv_whitebalance=%d" ADDCONFIG
			    description "��ƽ��: 1-Auto; 2-Fine; 3-Cloudy; 4-Filament Lamp; 5-Fluorescent Lamp"
		    }
		    
		    cdl_option dv_brightness {
			    display "brightness"
			    flavor data
			    no_define
			    default_value {"1"}
			    legal_values {"-3" "-2" "-1" "0" "1" "2" "3" }
			    define -format "dv_brightness=%d" ADDCONFIG
			    description "������: -3~3"
		    }
	    
		    cdl_option dv_exposure_mode {
			    display "exposure mode"
			    flavor data
			    no_define
			    default_value {"1"}
			    legal_values {"1" "2" "3"}
			    define -format "dv_exposure_mode=%d" ADDCONFIG
			    description "�ع�ģʽ: 1- Auto; 2-Indoor; 3-Outdoor"
		    }
		    
		    
		   
		    
        }
        
        cdl_component PC_CAMERA_CFG {
		    display "PC_CAMERA �������"
		    flavor none
		    no_define
		    description "PC_CAMERA���ѡ�������"
		
		    define_proc {
			    puts $::cdl_header ""
			    puts $::cdl_header "/*PC_CAMERA�������*/"
		    }
		    
        }
	    
	}
	
	cdl_component MUSIC_CFG {
		display "MUSIC �������"
		flavor none
		no_define
		description "MUSIC���ѡ�������"
		
		define_proc {
			puts $::cdl_header ""
			puts $::cdl_header "/*MUSIC�������*/"
		}
		
		cdl_option music_loop_mode {
			display "loop mode"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1" "2" "3" "4" "5"}
			define -format "music_loop_mode=%d" ADDCONFIG
			description "ѭ��ģʽ:0-Sequence, 1-Repeat All, 2-Repeat One, 3-Shuffle, 4-Shuffle + Repeat, 5-Intro"
		}
		
		cdl_option music_display_mode {
			display "display mode"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1" "2" "3" "4"}
			define -format "music_display_mode=%d" ADDCONFIG
			description "��ʾģʽ: 0-Spectrum, 1-Lyric, 2-Effect1, 3-Effect2, 4-Effect3"
		}
		
		cdl_option music_eq_mode {
			display "eq mode"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1" "2" "3" "4" "5" "6" "7" "8" "9" "10"}
			define -format "music_eq_mode=%d" ADDCONFIG
			description "Eq����:0-Norma, 1-Pop, 2-Classic, 3-Soft, 4-Jazz, 5-Rock, 6-DBB, 7-Custom EQ, 8-SRS WOW, 9-SRS WOW HD, 10-SRS USER Mode"
		}
		
		cdl_option music_srs_3d {
			display "srs 3d"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1" "2" "3" "4" "5" "6" "7" "8" "9" "10"}
			define -format "music_srs_3d=%d" ADDCONFIG
			description "Srs��srs 3dֵ:0 ~ 10"
		}
		
		cdl_option music_srs_trubass {
			display "srs trubass"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1" "2" "3" "4" "5" "6" "7" "8" "9" "10"}
			define -format "music_srs_trubass=%d" ADDCONFIG
			description "Srs��Trubassֵ:0 ~ 10"
		}
		
		cdl_option music_srs_focus {
			display "srs focus"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1" "2" "3" "4" "5" "6" "7" "8" "9" "10"}
			define -format "music_srs_focus=%d" ADDCONFIG
			description "Srs��Focusֵ:0 ~ 10"
		}
		
		cdl_option music_srs_center {
			display "srs center"
			flavor data
			no_define
			default_value {"1"}
			legal_values {"1" "2" "3" "4" "5" "6" "7" "8" "9" "10"}
			define -format "music_srs_center=%d" ADDCONFIG
			description "Srs��Centerֵ:1~ 10"
		}
		
		cdl_option music_srs_definition {
			display "srs definition"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1" "2" "3" "4" "5" "6" "7" "8" "9" "10"}
			define -format "music_srs_definition=%d" ADDCONFIG
			description "Srs��Definitionֵ:0 ~ 10"
		}
		
		cdl_option music_srs_speaker {
			display "srs speaker"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1" "2"}
			define -format "music_srs_speaker=%d" ADDCONFIG
			description "Srs��Speaker sizeֵ:0-60Hz, 1-100Hz, 2-150Hz"
		}
		
		cdl_option music_srs_limiter {
			display "srs limiter"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1"}
			define -format "music_srs_limiter=%d" ADDCONFIG
			description "Srs��Limiterֵ:0-disable, 1-enable"
		}
		
		cdl_option music_custom_80Hz {
			display "custom 80Hz"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"-6" "-5" "-4" "-3" "-2" "-1" "0" "1" "2" "3" "4" "5" "6"}
			define -format "music_custom_80Hz=%d" ADDCONFIG
			description "Custom Eq��80Hz����:-6db~+6db"
		}
		
		cdl_option music_custom_200Hz {
			display "custom 200Hz"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"-6" "-5" "-4" "-3" "-2" "-1" "0" "1" "2" "3" "4" "5" "6"}
			define -format "music_custom_200Hz=%d" ADDCONFIG
			description "Custom Eq��200Hz����:-6db~+6db"
		}
		
		cdl_option music_custom_1kHz {
			display "custom 1kHz"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"-6" "-5" "-4" "-3" "-2" "-1" "0" "1" "2" "3" "4" "5" "6"}
			define -format "music_custom_1kHz=%d" ADDCONFIG
			description "Custom Eq��1kHz����:-6db~+6db"
		}
		
		cdl_option music_custom_4kHz {
			display "custom 4kHz"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"-6" "-5" "-4" "-3" "-2" "-1" "0" "1" "2" "3" "4" "5" "6"}
			define -format "music_custom_4kHz=%d" ADDCONFIG
			description "Custom Eq��4kHz����:-6db~+6db"
		}
		
		cdl_option music_custom_8kHz {
			display "custom 8kHz"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"-6" "-5" "-4" "-3" "-2" "-1" "0" "1" "2" "3" "4" "5" "6"}
			define -format "music_custom_8kHz=%d" ADDCONFIG
			description "Custom Eq��8kHz����:-6db~+6db"
		}
		
		cdl_option music_fade {
			display "music fade"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1"}
			define -format "music_fade=%d" ADDCONFIG
			description "���뵭��:0-disable, 1-enable"
		}
		
		cdl_option music_speed {
			display "music speed"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"-4" "-3" "-2" "-1" "0" "1" "2" "3" "4"}
			define -format "music_speed=%d" ADDCONFIG
			description "���ٲ��ŵ��ٶ�:-4~+4"
		}
		
		cdl_option music_scan_speed {
			display "scan speed"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1" "2" "3" "4"}
			define -format "music_scan_speed=%d" ADDCONFIG
			description "ɨ���ٶ�:0-2X, 1-4X, 2-8X, 3-16X, 4-32X"
		}
		
	}
	
	cdl_component VIDEO_CFG {
		display "VIDEO �������"
		flavor none
		no_define
		description "VIDEO���ѡ�������"
		
		define_proc {
			puts $::cdl_header ""
			puts $::cdl_header "/*VIDEO�������*/"
		}
		
	}
	
	cdl_component EBOOK_CFG {
		display "EBOOK �������"
		flavor none
		no_define
		description "EBOOK���ѡ�������"
		
		define_proc {
			puts $::cdl_header ""
			puts $::cdl_header "/*EBOOK�������*/"
		}
		
		cdl_option ebook_roll_effect {
			display "roll effect"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1" "2"}
			define -format "ebook_roll_effect=%d" ADDCONFIG
			description "�Զ���������Ч: 0-�رգ�1-ƽ���Ϸ���2-���������ҳ"
		}
		
		cdl_option ebook_font_size {
			display "font size"
			flavor data
			no_define
			default_value {"12"}
			legal_values {"12" "16" "24"}
			define -format "ebook_font_size=%d" ADDCONFIG
			description "����Ĵ�С: 12-С��16-�У�24-��"
		}
		
		cdl_option ebook_font_color {
			display "font color"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1" "2" "3"}
			define -format "ebook_font_color=%d" ADDCONFIG
			description "�������ɫ: 0-���ף�1-��ɫ��2-���ң�3-����"
		}
	}
	
	cdl_component RECORD_CFG {
		display "RECORD �������"
		flavor none
		no_define
		description "RECORD���ѡ�������"
		
		define_proc {
			puts $::cdl_header ""
			puts $::cdl_header "/*RECORD�������*/"
		}
		
		cdl_option record_rectype {
			display "file type"
			flavor data
			no_define
			default_value {"0"}
			legal_values {"0" "1"}
			define -format "record_rectype=%d" ADDCONFIG
			description "¼���ļ���������: 0-wav;1-mp3"
		}
		
		cdl_option record_channel {
			display "channel"
			flavor data
			no_define
			default_value {"2"}
			legal_values {"1" "2"}
			define -format "record_channel=%d" ADDCONFIG
			description "��Ƶ������ͨ����:1-��������2-˫����"
		}
	}
	
	cdl_component TOOLS_CFG {
		display "TOOLS �������"
		flavor none
		no_define
		description "TOOLS���ѡ�������"
		
		define_proc {
			puts $::cdl_header ""
			puts $::cdl_header "/*TOOLS�������*/"
		}
		
		cdl_component CALENDAR_CFG {
		    display "CALENDAR �������"
		    flavor none
		    no_define
		    description "CALENDAR���ѡ�������"
		
		    define_proc {
			    puts $::cdl_header ""
			    puts $::cdl_header "/*CALENDAR�������*/"
		    }
		}	
		
		cdl_component STOPWATCH_CFG {
		    display "STOPWATCH �������"
		    flavor none
		    no_define
		    description "STOPWATCH���ѡ�������"
		
		    define_proc {
			    puts $::cdl_header ""
			    puts $::cdl_header "/*STOPWATCH�������*/"
		    }
		}	
		
		cdl_component CALCULATOR_CFG {
		    display "CALCULATOR �������"
		    flavor none
		    no_define
		    description "CALCULATOR���ѡ�������"
		
		    define_proc {
			    puts $::cdl_header ""
			    puts $::cdl_header "/*CALCULATOR�������*/"
		    }
		}	
		
	}
	
	cdl_component GAMES_CFG {
		display "GAMES �������"
		flavor none
		no_define
		description "GAMES���ѡ�������"
		
		define_proc {
			puts $::cdl_header ""
			puts $::cdl_header "/*GAMES�������*/"
		}
		cdl_component EMULATOR_CFG {
		    display "EMULATOR �������"
		    flavor none
		    no_define
		    description "EMULATOR���ѡ�������"
		
		    define_proc {
			    puts $::cdl_header ""
			    puts $::cdl_header "/*EMULATOR�������*/"
		    }
		}
		
		cdl_component G_GAME_CFG {
		    display "G_GAME �������"
		    flavor none
		    no_define
		    description "G_GAME���ѡ�������"
		
		    define_proc {
			    puts $::cdl_header ""
			    puts $::cdl_header "/*G_GAME�������*/"
		    }
		}	
		
	}
	
	cdl_component APPOTHERS_CFG {
		display "Ӧ�������������"
		flavor none
		no_define
		description "Ӧ���������ѡ�������"
		
		define_proc {
			puts $::cdl_header ""
			puts $::cdl_header "/*Ӧ�������������*/"
		}
		
	}
}

